magic
tech sky130A
magscale 1 2
timestamp 1727438411
<< viali >>
rect 3500 -630 4880 -590
rect 2430 -700 2590 -660
rect 2430 -2070 2590 -2030
rect 3500 -2070 4880 -2030
<< metal1 >>
rect 1800 -281 5800 -140
rect 1800 -380 5170 -281
rect 5269 -380 5800 -281
rect 1800 -460 5800 -380
rect 2110 -790 2240 -460
rect 2420 -640 2620 -460
rect 3150 -590 5130 -460
rect 3150 -630 3500 -590
rect 4880 -630 5130 -590
rect 3150 -640 5130 -630
rect 2410 -660 2630 -640
rect 2410 -700 2430 -660
rect 2590 -700 2630 -660
rect 2940 -700 5110 -690
rect 2410 -720 2630 -700
rect 2820 -740 5110 -700
rect 2110 -960 2490 -790
rect 2820 -800 2970 -740
rect 2540 -950 2970 -800
rect 3127 -842 3137 -787
rect 3193 -842 3203 -787
rect 3319 -842 3329 -787
rect 3385 -842 3395 -787
rect 3511 -842 3521 -787
rect 3577 -842 3587 -787
rect 3703 -842 3713 -787
rect 3769 -842 3779 -787
rect 3895 -842 3905 -787
rect 3961 -842 3971 -787
rect 4087 -842 4097 -787
rect 4153 -842 4163 -787
rect 4279 -842 4289 -787
rect 4345 -842 4355 -787
rect 4471 -842 4481 -787
rect 4537 -842 4547 -787
rect 4663 -842 4673 -787
rect 4729 -842 4739 -787
rect 4855 -842 4865 -787
rect 4921 -842 4931 -787
rect 5047 -844 5057 -789
rect 5119 -844 5129 -789
rect 2720 -1020 2970 -950
rect 3224 -956 3234 -900
rect 3295 -956 3305 -900
rect 3416 -956 3426 -900
rect 3487 -956 3497 -900
rect 3608 -956 3618 -900
rect 3679 -956 3689 -900
rect 3800 -956 3810 -900
rect 3871 -956 3881 -900
rect 3992 -956 4002 -900
rect 4063 -956 4073 -900
rect 4184 -956 4194 -900
rect 4255 -956 4265 -900
rect 4376 -956 4386 -900
rect 4447 -956 4457 -900
rect 4568 -956 4578 -900
rect 4639 -956 4649 -900
rect 4760 -956 4770 -900
rect 4831 -956 4841 -900
rect 4952 -956 4962 -900
rect 5023 -956 5033 -900
rect 2231 -1060 2539 -1021
rect 2231 -1200 2270 -1060
rect 1800 -1400 2270 -1200
rect 2231 -1680 2270 -1400
rect 2720 -1070 5110 -1020
rect 2720 -1610 2970 -1070
rect 5294 -1400 5300 -1200
rect 5500 -1400 5800 -1200
rect 2720 -1660 5110 -1610
rect 2231 -1719 2539 -1680
rect 2160 -1910 2490 -1770
rect 2720 -1780 2970 -1660
rect 3124 -1761 3134 -1706
rect 3190 -1761 3200 -1706
rect 3316 -1761 3326 -1706
rect 3382 -1761 3392 -1706
rect 3508 -1761 3518 -1706
rect 3574 -1761 3584 -1706
rect 3700 -1761 3710 -1706
rect 3766 -1761 3776 -1706
rect 3892 -1761 3902 -1706
rect 3958 -1761 3968 -1706
rect 4084 -1761 4094 -1706
rect 4150 -1761 4160 -1706
rect 4276 -1761 4286 -1706
rect 4342 -1761 4352 -1706
rect 4468 -1761 4478 -1706
rect 4534 -1761 4544 -1706
rect 4660 -1761 4670 -1706
rect 4726 -1761 4736 -1706
rect 4852 -1761 4862 -1706
rect 4918 -1761 4928 -1706
rect 5047 -1763 5057 -1708
rect 5119 -1763 5129 -1708
rect 2160 -2140 2300 -1910
rect 2530 -1920 2970 -1780
rect 3221 -1875 3231 -1819
rect 3292 -1875 3302 -1819
rect 3413 -1875 3423 -1819
rect 3484 -1875 3494 -1819
rect 3605 -1875 3615 -1819
rect 3676 -1875 3686 -1819
rect 3797 -1875 3807 -1819
rect 3868 -1875 3878 -1819
rect 3989 -1875 3999 -1819
rect 4060 -1875 4070 -1819
rect 4181 -1875 4191 -1819
rect 4252 -1875 4262 -1819
rect 4373 -1875 4383 -1819
rect 4444 -1875 4454 -1819
rect 4565 -1875 4575 -1819
rect 4636 -1875 4646 -1819
rect 4757 -1875 4767 -1819
rect 4828 -1875 4838 -1819
rect 4949 -1875 4959 -1819
rect 5020 -1875 5030 -1819
rect 2530 -1930 5110 -1920
rect 2820 -1970 5110 -1930
rect 2410 -2030 2620 -2010
rect 2410 -2070 2430 -2030
rect 2590 -2070 2620 -2030
rect 2420 -2140 2620 -2070
rect 3140 -2030 5120 -2020
rect 3140 -2070 3500 -2030
rect 4880 -2070 5120 -2030
rect 3140 -2140 5120 -2070
rect 1800 -2155 5800 -2140
rect 1800 -2305 5145 -2155
rect 5295 -2305 5800 -2155
rect 1800 -2460 5800 -2305
<< via1 >>
rect 5170 -380 5269 -281
rect 3137 -842 3193 -787
rect 3329 -842 3385 -787
rect 3521 -842 3577 -787
rect 3713 -842 3769 -787
rect 3905 -842 3961 -787
rect 4097 -842 4153 -787
rect 4289 -842 4345 -787
rect 4481 -842 4537 -787
rect 4673 -842 4729 -787
rect 4865 -842 4921 -787
rect 5057 -844 5119 -789
rect 3234 -956 3295 -900
rect 3426 -956 3487 -900
rect 3618 -956 3679 -900
rect 3810 -956 3871 -900
rect 4002 -956 4063 -900
rect 4194 -956 4255 -900
rect 4386 -956 4447 -900
rect 4578 -956 4639 -900
rect 4770 -956 4831 -900
rect 4962 -956 5023 -900
rect 5300 -1400 5500 -1200
rect 3134 -1761 3190 -1706
rect 3326 -1761 3382 -1706
rect 3518 -1761 3574 -1706
rect 3710 -1761 3766 -1706
rect 3902 -1761 3958 -1706
rect 4094 -1761 4150 -1706
rect 4286 -1761 4342 -1706
rect 4478 -1761 4534 -1706
rect 4670 -1761 4726 -1706
rect 4862 -1761 4918 -1706
rect 5057 -1763 5119 -1708
rect 3231 -1875 3292 -1819
rect 3423 -1875 3484 -1819
rect 3615 -1875 3676 -1819
rect 3807 -1875 3868 -1819
rect 3999 -1875 4060 -1819
rect 4191 -1875 4252 -1819
rect 4383 -1875 4444 -1819
rect 4575 -1875 4636 -1819
rect 4767 -1875 4828 -1819
rect 4959 -1875 5020 -1819
rect 5145 -2305 5295 -2155
<< metal2 >>
rect 5170 -281 5269 -275
rect 5170 -690 5269 -380
rect 3120 -787 5269 -690
rect 3120 -842 3137 -787
rect 3193 -842 3329 -787
rect 3385 -842 3521 -787
rect 3577 -842 3713 -787
rect 3769 -842 3905 -787
rect 3961 -842 4097 -787
rect 4153 -842 4289 -787
rect 4345 -842 4481 -787
rect 4537 -842 4673 -787
rect 4729 -842 4865 -787
rect 4921 -789 5269 -787
rect 4921 -842 5057 -789
rect 3120 -844 5057 -842
rect 5119 -844 5180 -789
rect 3120 -850 5180 -844
rect 3137 -852 3193 -850
rect 3329 -852 3385 -850
rect 3521 -852 3577 -850
rect 3713 -852 3769 -850
rect 3905 -852 3961 -850
rect 4097 -852 4153 -850
rect 4289 -852 4345 -850
rect 4481 -852 4537 -850
rect 4673 -852 4729 -850
rect 4865 -852 4921 -850
rect 5057 -854 5119 -850
rect 3120 -900 5174 -890
rect 3120 -956 3234 -900
rect 3295 -956 3426 -900
rect 3487 -956 3618 -900
rect 3679 -956 3810 -900
rect 3871 -956 4002 -900
rect 4063 -956 4194 -900
rect 4255 -956 4386 -900
rect 4447 -956 4578 -900
rect 4639 -956 4770 -900
rect 4831 -956 4962 -900
rect 5023 -956 5174 -900
rect 3120 -960 5174 -956
rect 3120 -1060 5170 -960
rect 5000 -1200 5170 -1060
rect 5300 -1200 5500 -1194
rect 5000 -1400 5300 -1200
rect 5000 -1580 5170 -1400
rect 5300 -1406 5500 -1400
rect 3120 -1699 5170 -1580
rect 3117 -1706 5171 -1699
rect 3117 -1761 3134 -1706
rect 3190 -1761 3326 -1706
rect 3382 -1761 3518 -1706
rect 3574 -1761 3710 -1706
rect 3766 -1761 3902 -1706
rect 3958 -1761 4094 -1706
rect 4150 -1761 4286 -1706
rect 4342 -1761 4478 -1706
rect 4534 -1761 4670 -1706
rect 4726 -1761 4862 -1706
rect 4918 -1708 5171 -1706
rect 4918 -1761 5057 -1708
rect 3117 -1763 5057 -1761
rect 5119 -1763 5171 -1708
rect 3117 -1769 5171 -1763
rect 3134 -1771 3190 -1769
rect 3326 -1771 3382 -1769
rect 3518 -1771 3574 -1769
rect 3710 -1771 3766 -1769
rect 3902 -1771 3958 -1769
rect 4094 -1771 4150 -1769
rect 4286 -1771 4342 -1769
rect 4478 -1771 4534 -1769
rect 4670 -1771 4726 -1769
rect 4862 -1771 4918 -1769
rect 5057 -1773 5119 -1769
rect 3117 -1819 5171 -1809
rect 3117 -1875 3231 -1819
rect 3292 -1875 3423 -1819
rect 3484 -1875 3615 -1819
rect 3676 -1875 3807 -1819
rect 3868 -1875 3999 -1819
rect 4060 -1875 4191 -1819
rect 4252 -1875 4383 -1819
rect 4444 -1875 4575 -1819
rect 4636 -1875 4767 -1819
rect 4828 -1875 4959 -1819
rect 5020 -1830 5171 -1819
rect 5020 -1875 5295 -1830
rect 3117 -1879 5295 -1875
rect 3120 -1980 5295 -1879
rect 5145 -2155 5295 -1980
rect 5145 -2311 5295 -2305
use sky130_fd_pr__pfet_01v8_2DVCWQ  sky130_fd_pr__pfet_01v8_2DVCWQ_0
timestamp 1727436632
transform 1 0 4127 0 1 -881
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_MGS3BN  XM1
timestamp 1727436632
transform 1 0 2511 0 -1 -916
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1727436632
transform 1 0 2511 0 1 -1821
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_FUP3AZ  XM4
timestamp 1727438070
transform 1 0 4127 0 1 -1790
box -1127 -310 1127 310
<< labels >>
flabel metal1 5600 -1400 5800 -1200 0 FreeSans 256 0 0 0 output
port 2 nsew
flabel metal1 1800 -1400 2000 -1200 0 FreeSans 256 0 0 0 input
port 3 nsew
flabel metal1 1860 -380 2060 -180 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1860 -2380 2060 -2180 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 2720 -1890 2840 -830 0 FreeSans 320 0 0 0 inverted
<< end >>
